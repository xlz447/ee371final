library verilog;
use verilog.vl_types.all;
entity clkCounter_vlg_vec_tst is
end clkCounter_vlg_vec_tst;
