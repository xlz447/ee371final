library verilog;
use verilog.vl_types.all;
entity clkCounter2_vlg_vec_tst is
end clkCounter2_vlg_vec_tst;
